module top_module (
    input clk, d,
    output q);

    

endmodule