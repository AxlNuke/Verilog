module top_module ( input a, input b, output out );
    mod_a instancia1 (a, b, out);
endmodule